`ifndef _PARAMS_VH_
`define _PARAMS_VH_

// game state
parameter GS_INIT         = 4'd0;
parameter GS_IDLE         = 4'd1;
parameter GS_RELOAD       = 4'd2;

parameter TILE_BLANK      = 8'd0;
parameter TILE_WALL       = 8'd1;

`endif