`ifndef _PARAMS_VH_
`define _PARAMS_VH_

parameter TILE_BLANK      = 8'd0;
parameter TILE_WALL       = 8'd1;



`endif