
module CLK_25M (
	clk_clk,
	reset_reset_n,
	clk_25m_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		clk_25m_clk;
endmodule
